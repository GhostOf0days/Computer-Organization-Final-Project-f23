`timescale 1 ns / 1 ps

module test_cpu;
    parameter 